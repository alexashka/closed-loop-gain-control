/*
  sync_rom  rom_label(
    .clk(clk), 
	.address(), 
	.data_out());
*/
module sync_rom(clk, address, data_out);
  input clk;
  input [7:0] address;
  output [7:0] data_out;
  // local ///
  reg [7:0] data_out;
  always @ (posedge clk) begin
    case (address)
    8'b0: data_out <= 8'b1;
    8'b1: data_out <= 8'b10;
    8'b10: data_out <= 8'b100;
    8'b11: data_out <= 8'b1000;
    8'b100: data_out <= 8'b10000;
    8'b101: data_out <= 8'b100000;
    8'b110: data_out <= 8'b1000000;
    8'b111: data_out <= 8'b10000000;
    8'b1000: data_out <= 8'b11101;
    8'b1001: data_out <= 8'b111010;
    8'b1010: data_out <= 8'b1110100;
    8'b1011: data_out <= 8'b11101000;
    8'b1100: data_out <= 8'b11001101;
    8'b1101: data_out <= 8'b10000111;
    8'b1110: data_out <= 8'b10011;
    8'b1111: data_out <= 8'b100110;
    8'b10000: data_out <= 8'b1001100;
    8'b10001: data_out <= 8'b10011000;
    8'b10010: data_out <= 8'b101101;
    8'b10011: data_out <= 8'b1011010;
    8'b10100: data_out <= 8'b10110100;
    8'b10101: data_out <= 8'b1110101;
    8'b10110: data_out <= 8'b11101010;
    8'b10111: data_out <= 8'b11001001;
    8'b11000: data_out <= 8'b10001111;
    8'b11001: data_out <= 8'b11;
    8'b11010: data_out <= 8'b110;
    8'b11011: data_out <= 8'b1100;
    8'b11100: data_out <= 8'b11000;
    8'b11101: data_out <= 8'b110000;
    8'b11110: data_out <= 8'b1100000;
    8'b11111: data_out <= 8'b11000000;
    8'b100000: data_out <= 8'b10011101;
    8'b100001: data_out <= 8'b100111;
    8'b100010: data_out <= 8'b1001110;
    8'b100011: data_out <= 8'b10011100;
    8'b100100: data_out <= 8'b100101;
    8'b100101: data_out <= 8'b1001010;
    8'b100110: data_out <= 8'b10010100;
    8'b100111: data_out <= 8'b110101;
    8'b101000: data_out <= 8'b1101010;
    8'b101001: data_out <= 8'b11010100;
    8'b101010: data_out <= 8'b10110101;
    8'b101011: data_out <= 8'b1110111;
    8'b101100: data_out <= 8'b11101110;
    8'b101101: data_out <= 8'b11000001;
    8'b101110: data_out <= 8'b10011111;
    8'b101111: data_out <= 8'b100011;
    8'b110000: data_out <= 8'b1000110;
    8'b110001: data_out <= 8'b10001100;
    8'b110010: data_out <= 8'b101;
    8'b110011: data_out <= 8'b1010;
    8'b110100: data_out <= 8'b10100;
    8'b110101: data_out <= 8'b101000;
    8'b110110: data_out <= 8'b1010000;
    8'b110111: data_out <= 8'b10100000;
    8'b111000: data_out <= 8'b1011101;
    8'b111001: data_out <= 8'b10111010;
    8'b111010: data_out <= 8'b1101001;
    8'b111011: data_out <= 8'b11010010;
    8'b111100: data_out <= 8'b10111001;
    8'b111101: data_out <= 8'b1101111;
    8'b111110: data_out <= 8'b11011110;
    8'b111111: data_out <= 8'b10100001;
    8'b1000000: data_out <= 8'b1011111;
    8'b1000001: data_out <= 8'b10111110;
    8'b1000010: data_out <= 8'b1100001;
    8'b1000011: data_out <= 8'b11000010;
    8'b1000100: data_out <= 8'b10011001;
    8'b1000101: data_out <= 8'b101111;
    8'b1000110: data_out <= 8'b1011110;
    8'b1000111: data_out <= 8'b10111100;
    8'b1001000: data_out <= 8'b1100101;
    8'b1001001: data_out <= 8'b11001010;
    8'b1001010: data_out <= 8'b10001001;
    8'b1001011: data_out <= 8'b1111;
    8'b1001100: data_out <= 8'b11110;
    8'b1001101: data_out <= 8'b111100;
    8'b1001110: data_out <= 8'b1111000;
    8'b1001111: data_out <= 8'b11110000;
    8'b1010000: data_out <= 8'b11111101;
    8'b1010001: data_out <= 8'b11100111;
    8'b1010010: data_out <= 8'b11010011;
    8'b1010011: data_out <= 8'b10111011;
    8'b1010100: data_out <= 8'b1101011;
    8'b1010101: data_out <= 8'b11010110;
    8'b1010110: data_out <= 8'b10110001;
    8'b1010111: data_out <= 8'b1111111;
    8'b1011000: data_out <= 8'b11111110;
    8'b1011001: data_out <= 8'b11100001;
    8'b1011010: data_out <= 8'b11011111;
    8'b1011011: data_out <= 8'b10100011;
    8'b1011100: data_out <= 8'b1011011;
    8'b1011101: data_out <= 8'b10110110;
    8'b1011110: data_out <= 8'b1110001;
    8'b1011111: data_out <= 8'b11100010;
    8'b1100000: data_out <= 8'b11011001;
    8'b1100001: data_out <= 8'b10101111;
    8'b1100010: data_out <= 8'b1000011;
    8'b1100011: data_out <= 8'b10000110;
    8'b1100100: data_out <= 8'b10001;
    8'b1100101: data_out <= 8'b100010;
    8'b1100110: data_out <= 8'b1000100;
    8'b1100111: data_out <= 8'b10001000;
    8'b1101000: data_out <= 8'b1101;
    8'b1101001: data_out <= 8'b11010;
    8'b1101010: data_out <= 8'b110100;
    8'b1101011: data_out <= 8'b1101000;
    8'b1101100: data_out <= 8'b11010000;
    8'b1101101: data_out <= 8'b10111101;
    8'b1101110: data_out <= 8'b1100111;
    8'b1101111: data_out <= 8'b11001110;
    8'b1110000: data_out <= 8'b10000001;
    8'b1110001: data_out <= 8'b11111;
    8'b1110010: data_out <= 8'b111110;
    8'b1110011: data_out <= 8'b1111100;
    8'b1110100: data_out <= 8'b11111000;
    8'b1110101: data_out <= 8'b11101101;
    8'b1110110: data_out <= 8'b11000111;
    8'b1110111: data_out <= 8'b10010011;
    8'b1111000: data_out <= 8'b111011;
    8'b1111001: data_out <= 8'b1110110;
    8'b1111010: data_out <= 8'b11101100;
    8'b1111011: data_out <= 8'b11000101;
    8'b1111100: data_out <= 8'b10010111;
    8'b1111101: data_out <= 8'b110011;
    8'b1111110: data_out <= 8'b1100110;
    8'b1111111: data_out <= 8'b11001100;
    8'b10000000: data_out <= 8'b10000101;
    8'b10000001: data_out <= 8'b10111;
    8'b10000010: data_out <= 8'b101110;
    8'b10000011: data_out <= 8'b1011100;
    8'b10000100: data_out <= 8'b10111000;
    8'b10000101: data_out <= 8'b1101101;
    8'b10000110: data_out <= 8'b11011010;
    8'b10000111: data_out <= 8'b10101001;
    8'b10001000: data_out <= 8'b1001111;
    8'b10001001: data_out <= 8'b10011110;
    8'b10001010: data_out <= 8'b100001;
    8'b10001011: data_out <= 8'b1000010;
    8'b10001100: data_out <= 8'b10000100;
    8'b10001101: data_out <= 8'b10101;
    8'b10001110: data_out <= 8'b101010;
    8'b10001111: data_out <= 8'b1010100;
    8'b10010000: data_out <= 8'b10101000;
    8'b10010001: data_out <= 8'b1001101;
    8'b10010010: data_out <= 8'b10011010;
    8'b10010011: data_out <= 8'b101001;
    8'b10010100: data_out <= 8'b1010010;
    8'b10010101: data_out <= 8'b10100100;
    8'b10010110: data_out <= 8'b1010101;
    8'b10010111: data_out <= 8'b10101010;
    8'b10011000: data_out <= 8'b1001001;
    8'b10011001: data_out <= 8'b10010010;
    8'b10011010: data_out <= 8'b111001;
    8'b10011011: data_out <= 8'b1110010;
    8'b10011100: data_out <= 8'b11100100;
    8'b10011101: data_out <= 8'b11010101;
    8'b10011110: data_out <= 8'b10110111;
    8'b10011111: data_out <= 8'b1110011;
    8'b10100000: data_out <= 8'b11100110;
    8'b10100001: data_out <= 8'b11010001;
    8'b10100010: data_out <= 8'b10111111;
    8'b10100011: data_out <= 8'b1100011;
    8'b10100100: data_out <= 8'b11000110;
    8'b10100101: data_out <= 8'b10010001;
    8'b10100110: data_out <= 8'b111111;
    8'b10100111: data_out <= 8'b1111110;
    8'b10101000: data_out <= 8'b11111100;
    8'b10101001: data_out <= 8'b11100101;
    8'b10101010: data_out <= 8'b11010111;
    8'b10101011: data_out <= 8'b10110011;
    8'b10101100: data_out <= 8'b1111011;
    8'b10101101: data_out <= 8'b11110110;
    8'b10101110: data_out <= 8'b11110001;
    8'b10101111: data_out <= 8'b11111111;
    8'b10110000: data_out <= 8'b11100011;
    8'b10110001: data_out <= 8'b11011011;
    8'b10110010: data_out <= 8'b10101011;
    8'b10110011: data_out <= 8'b1001011;
    8'b10110100: data_out <= 8'b10010110;
    8'b10110101: data_out <= 8'b110001;
    8'b10110110: data_out <= 8'b1100010;
    8'b10110111: data_out <= 8'b11000100;
    8'b10111000: data_out <= 8'b10010101;
    8'b10111001: data_out <= 8'b110111;
    8'b10111010: data_out <= 8'b1101110;
    8'b10111011: data_out <= 8'b11011100;
    8'b10111100: data_out <= 8'b10100101;
    8'b10111101: data_out <= 8'b1010111;
    8'b10111110: data_out <= 8'b10101110;
    8'b10111111: data_out <= 8'b1000001;
    8'b11000000: data_out <= 8'b10000010;
    8'b11000001: data_out <= 8'b11001;
    8'b11000010: data_out <= 8'b110010;
    8'b11000011: data_out <= 8'b1100100;
    8'b11000100: data_out <= 8'b11001000;
    8'b11000101: data_out <= 8'b10001101;
    8'b11000110: data_out <= 8'b111;
    8'b11000111: data_out <= 8'b1110;
    8'b11001000: data_out <= 8'b11100;
    8'b11001001: data_out <= 8'b111000;
    8'b11001010: data_out <= 8'b1110000;
    8'b11001011: data_out <= 8'b11100000;
    8'b11001100: data_out <= 8'b11011101;
    8'b11001101: data_out <= 8'b10100111;
    8'b11001110: data_out <= 8'b1010011;
    8'b11001111: data_out <= 8'b10100110;
    8'b11010000: data_out <= 8'b1010001;
    8'b11010001: data_out <= 8'b10100010;
    8'b11010010: data_out <= 8'b1011001;
    8'b11010011: data_out <= 8'b10110010;
    8'b11010100: data_out <= 8'b1111001;
    8'b11010101: data_out <= 8'b11110010;
    8'b11010110: data_out <= 8'b11111001;
    8'b11010111: data_out <= 8'b11101111;
    8'b11011000: data_out <= 8'b11000011;
    8'b11011001: data_out <= 8'b10011011;
    8'b11011010: data_out <= 8'b101011;
    8'b11011011: data_out <= 8'b1010110;
    8'b11011100: data_out <= 8'b10101100;
    8'b11011101: data_out <= 8'b1000101;
    8'b11011110: data_out <= 8'b10001010;
    8'b11011111: data_out <= 8'b1001;
    8'b11100000: data_out <= 8'b10010;
    8'b11100001: data_out <= 8'b100100;
    8'b11100010: data_out <= 8'b1001000;
    8'b11100011: data_out <= 8'b10010000;
    8'b11100100: data_out <= 8'b111101;
    8'b11100101: data_out <= 8'b1111010;
    8'b11100110: data_out <= 8'b11110100;
    8'b11100111: data_out <= 8'b11110101;
    8'b11101000: data_out <= 8'b11110111;
    8'b11101001: data_out <= 8'b11110011;
    8'b11101010: data_out <= 8'b11111011;
    8'b11101011: data_out <= 8'b11101011;
    8'b11101100: data_out <= 8'b11001011;
    8'b11101101: data_out <= 8'b10001011;
    8'b11101110: data_out <= 8'b1011;
    8'b11101111: data_out <= 8'b10110;
    8'b11110000: data_out <= 8'b101100;
    8'b11110001: data_out <= 8'b1011000;
    8'b11110010: data_out <= 8'b10110000;
    8'b11110011: data_out <= 8'b1111101;
    8'b11110100: data_out <= 8'b11111010;
    8'b11110101: data_out <= 8'b11101001;
    8'b11110110: data_out <= 8'b11001111;
    8'b11110111: data_out <= 8'b10000011;
    8'b11111000: data_out <= 8'b11011;
    8'b11111001: data_out <= 8'b110110;
    8'b11111010: data_out <= 8'b1101100;
    8'b11111011: data_out <= 8'b11011000;
    8'b11111100: data_out <= 8'b10101101;
    8'b11111101: data_out <= 8'b1000111;
    8'b11111110: data_out <= 8'b10001110;
    8'b11111111: data_out <= 8'b0;
    endcase
  end
endmodule
